* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_4 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.0707237516550235u tpotv=2.135726333967107n tpwv=230.47701920458005n 
    + tnln=0.0714282663367119u tnwn=139.8358833754729n tnotv=1.7293994430296098n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06093749048307959u tpotv=1.9903188745659293n tpwv=222.45071662992666n 
    + tnln=0.06179674979765479u tnwn=145.6270098559658n tnotv=1.6990599927247585n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06933208142952162u tpotv=2.062021322689429n tpwv=230.1089247173208n 
    + tnln=0.061071209277942386u tnwn=110.89677990857533n tnotv=1.941036078244934n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06993619034409022u tpotv=1.915720328710461n tpwv=236.61436687592334n 
    + tnln=0.062419869772087466u tnwn=118.25561325247398n tnotv=1.82993056296588n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.063857062413318u tpotv=1.763058478552256n tpwv=233.40468395492343n 
    + tnln=0.06108512235403309u tnwn=146.6304513732537n tnotv=1.7603593766832524n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.07060359066871835u tpotv=2.138638840144838n tpwv=237.9715498506643n 
    + tnln=0.07268608768452992u tnwn=119.64770639660824n tnotv=2.012628828583122n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06967049955850103u tpotv=2.048766518823419n tpwv=240.1552169178878n 
    + tnln=0.06658412747664814u tnwn=121.18430643048103n tnotv=1.8155698967172165n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.05552430302187232u tpotv=1.9710974037041011n tpwv=243.8724084313829n 
    + tnln=0.07305900253943082u tnwn=132.94067387096652n tnotv=1.7671486398478151n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.05564398065589843u tpotv=1.8246254311923988n tpwv=191.73674710190204n 
    + tnln=0.055515629660465526u tnwn=110.55574353484221n tnotv=1.844002139261351n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06761774297112173u tpotv=1.8411637046735891n tpwv=218.99158293114604n 
    + tnln=0.06428891454429068u tnwn=119.87458689088766n tnotv=1.9158560981740653n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.05972971073055329u tpotv=1.8053637862340748n tpwv=250.55025678547165n 
    + tnln=0.06327963035210127u tnwn=130.1969243323308n tnotv=1.7380610467900959n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.0740876723876319u tpotv=2.0625925427726752n tpwv=190.96865613461995n 
    + tnln=0.07017571865478416u tnwn=144.85367768283837n tnotv=1.7867401446741042n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.057897278523802005u tpotv=2.050961043231565n tpwv=235.3662932575614n 
    + tnln=0.060850798721719376u tnwn=138.23798768608108n tnotv=2.0144451101643974n 

.ENDS ring_osc.end
