* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_6 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.07414606444039876u tpotv=2.049098285027006n tpwv=233.6472557450415n 
    + tnln=0.07204441639064935u tnwn=140.42464359851962n tnotv=1.9115201798437296n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.07364113523180521u tpotv=2.1301051649534357n tpwv=207.66038704830362n 
    + tnln=0.07009547708429502u tnwn=125.85815171920245n tnotv=1.7393593222204329n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06574292629426495u tpotv=2.0858610222236758n tpwv=186.22047257278666n 
    + tnln=0.055323230523873376u tnwn=135.6196677154246n tnotv=1.9508716235336814n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06950092101006014u tpotv=2.1111844448474515n tpwv=241.5529002114007n 
    + tnln=0.06839605458300034u tnwn=126.1181818748841n tnotv=1.916178345314334n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.062184852120937176u tpotv=2.05596150323273n tpwv=208.3976574902857n 
    + tnln=0.06744907973343028u tnwn=147.72835625606976n tnotv=1.8148959135007012n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.05708920417655955u tpotv=1.890484792147543n tpwv=242.35678026188987n 
    + tnln=0.05682618458551668u tnwn=126.19880214097235n tnotv=1.679898653942641n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.0694555841505055u tpotv=1.9800578168227478n tpwv=212.2257502927167n 
    + tnln=0.059080549847877147u tnwn=138.2205658414459n tnotv=1.99939603796091n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.07004004588832644u tpotv=1.9850055688453943n tpwv=196.53702251493524n 
    + tnln=0.060741289013456795u tnwn=136.49295869712972n tnotv=1.7907359718273488n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.0679787843803653u tpotv=1.9747315489404924n tpwv=194.9796706997053n 
    + tnln=0.06215164225185987u tnwn=121.03975840372459n tnotv=1.9386069497290341n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.05578392587361866u tpotv=2.1424281494080946n tpwv=208.07965760963717n 
    + tnln=0.07047430706727993u tnwn=110.67015395710094n tnotv=1.8586349693891002n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.05865341079202198u tpotv=1.9336092584065803n tpwv=242.0486703546783n 
    + tnln=0.05847655271033048u tnwn=117.58542698890946n tnotv=1.8254232335235683n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.06302285195295208u tpotv=1.8865520987155224n tpwv=199.95298902419145n 
    + tnln=0.0705033865207119u tnwn=148.63374983368018n tnotv=1.9769293293215413n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06044215958981158u tpotv=1.8748303429936062n tpwv=218.88982273140562n 
    + tnln=0.07015170435665728u tnwn=125.01630924222883n tnotv=1.977505989403657n 

.ENDS ring_osc.end
