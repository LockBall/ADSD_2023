* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_1 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.06603835361641834u tpotv=1.8861382963862796n tpwv=204.39342127438061n 
    + tnln=0.0648194955662437u tnwn=132.28235674144096n tnotv=1.8812600980220011n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06327875845576124u tpotv=1.9312076948132189n tpwv=224.77223894518966n 
    + tnln=0.06189974288430767u tnwn=123.35689513383022n tnotv=1.666912720603328n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.0603251495489811u tpotv=1.8597764306276372n tpwv=223.4745756982782n 
    + tnln=0.07233673132349683u tnwn=126.93981414230176n tnotv=1.8991831590164914n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.05979343373236621u tpotv=1.7572183266005639n tpwv=202.69783278842164n 
    + tnln=0.05847926675074214u tnwn=121.81349596490584n tnotv=1.7693186562031449n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.06256844908587786u tpotv=1.764564749191225n tpwv=219.72588564617234n 
    + tnln=0.06120799007760081u tnwn=132.60048172371893n tnotv=1.9245960761437875n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06909909949145741u tpotv=1.856391304772322n tpwv=213.61884842986407n 
    + tnln=0.055387009520374286u tnwn=139.4191890594769n tnotv=1.9732985077591136n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.05875872566783576u tpotv=2.0530200667829974n tpwv=235.20806681483705n 
    + tnln=0.06994037844074655u tnwn=144.31058053916885n tnotv=1.736248547188473n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06517615576267774u tpotv=1.8471655782636895n tpwv=246.815536765962n 
    + tnln=0.06938751862243338u tnwn=139.43833567022523n tnotv=1.6796738761268446n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06088457774307084u tpotv=1.8562475757146653n tpwv=214.31588726855696n 
    + tnln=0.07402794183507627u tnwn=132.4520242188418n tnotv=1.6879056488906432n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06617323170766967u tpotv=1.9832019994908041n tpwv=225.2388367068748n 
    + tnln=0.05803210848118025u tnwn=131.07680927863328n tnotv=1.7866261769639622n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06207489998667842u tpotv=2.136518443802609n tpwv=245.8688457707903n 
    + tnln=0.07445356083881866u tnwn=123.41357855416743n tnotv=1.9920056340501355n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.05586621215038255u tpotv=1.948726835491152n tpwv=206.65531189398695n 
    + tnln=0.06959726795807568u tnwn=145.4314685975n tnotv=1.926846429563997n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.05911227616706696u tpotv=1.826702144835872n tpwv=205.94795743998682n 
    + tnln=0.06662682377508151u tnwn=123.79128002695333n tnotv=1.7361178359749183n 

.ENDS ring_osc.end
