* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_2 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.05609165919482345u tpotv=1.8653895105989944n tpwv=249.03495787711543n 
    + tnln=0.05940540629790855u tnwn=149.10004220471168n tnotv=1.99800703286893n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06045901844753077u tpotv=1.9949502112951278n tpwv=185.975956794318n 
    + tnln=0.05956421587110726u tnwn=133.58154941952574n tnotv=1.9065315777825675n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06251111025492083u tpotv=1.921193321183554n tpwv=219.38560702594592n 
    + tnln=0.06563108222983387u tnwn=116.49410630717921n tnotv=1.880214652645602n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.07457377419886255u tpotv=1.8038967285315526n tpwv=209.42215273712424n 
    + tnln=0.07283917057201864u tnwn=125.91149211918643n tnotv=1.94778228538215n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.065194665337686u tpotv=1.869269436508786n tpwv=242.27301099125668n 
    + tnln=0.06953446053305447u tnwn=120.20622491642851n tnotv=1.8033360099032614n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06067979703789237u tpotv=2.112177913680706n tpwv=216.5390324277805n 
    + tnln=0.071755459172121u tnwn=133.67263068165022n tnotv=1.7999474311910773n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06457771395984895u tpotv=1.800620025755232n tpwv=190.08836226443432n 
    + tnln=0.0600200106983982u tnwn=129.08604206641027n tnotv=1.767122094426043n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06861605354066194u tpotv=1.882742479595101n tpwv=224.5348924396552n 
    + tnln=0.05717759600306395u tnwn=145.93544162235932n tnotv=1.7844812466075566n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06747902599380291u tpotv=2.021061514435238n tpwv=190.5738965586211n 
    + tnln=0.0707730278611958u tnwn=112.67959639006835n tnotv=1.781929608344992n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.05593456779371392u tpotv=1.8520861004920952n tpwv=186.74083985537675n 
    + tnln=0.07022442989549894u tnwn=128.54681610534794n tnotv=1.9931983101701225n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06765552921723411u tpotv=2.0238458995713473n tpwv=223.89597137992504n 
    + tnln=0.06036416750558327u tnwn=118.31729370715998n tnotv=1.6727394624657717n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.05685595411638272u tpotv=1.9699095774840767n tpwv=235.54829395545877n 
    + tnln=0.06719744949139608u tnwn=115.51717429636113n tnotv=1.7623939410403193n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06878142025033365u tpotv=2.102751523452824n tpwv=247.46187751622588n 
    + tnln=0.07251141534594435u tnwn=135.97478603374395n tnotv=1.6766425782739591n 

.ENDS ring_osc.end
