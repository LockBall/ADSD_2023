library ieee;
use ieee.std_logic_1164.all;

entity proj_5 is

    port(
        clk: in std_logic;
        reset_n: std_logic
    );

end entity;


architecture arch of proj_5 is



begin
end architecture;