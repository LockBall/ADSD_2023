* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_3 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.055959387641422983u tpotv=1.7571902371251937n tpwv=188.7144203533245n 
    + tnln=0.0572434841139237u tnwn=120.30175336370678n tnotv=1.9808170892044312n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.07455329653432445u tpotv=2.009534646497045n tpwv=240.02361431066274n 
    + tnln=0.07177783261062928u tnwn=146.04576494638482n tnotv=1.683986415863397n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06708932728008564u tpotv=1.8045142998056996n tpwv=212.3180503575455n 
    + tnln=0.05605666109840014u tnwn=134.55825452710516n tnotv=1.791972982566331n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.059350863799019674u tpotv=1.8843059378151283n tpwv=202.68374429631922n 
    + tnln=0.06699691107050862u tnwn=138.274230643894n tnotv=2.0170043715596617n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.06195655183453155u tpotv=1.9984084336584333n tpwv=238.1386358440064n 
    + tnln=0.07077612514964789u tnwn=119.10505493810946n tnotv=1.8540597940558627n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06116115969119908u tpotv=1.7589068521534823n tpwv=211.04057057323985n 
    + tnln=0.06240440114368234u tnwn=119.45554943575252n tnotv=1.8824890897591882n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06932476618955394u tpotv=1.9491880888840754n tpwv=200.12724025962603n 
    + tnln=0.0741461525953223u tnwn=147.09416958952096n tnotv=1.981929895796839n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06622200560052009u tpotv=2.0929717441818574n tpwv=201.2952218722724n 
    + tnln=0.06919765213945264u tnwn=124.74212823429927n tnotv=1.8906703265498364n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.0680592884526949u tpotv=2.139437268970906n tpwv=185.983114195254n 
    + tnln=0.0569157705295487u tnwn=114.48567839032462n tnotv=1.9018273362196312n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0672042766393191u tpotv=2.0158369887317042n tpwv=246.54542027989524n 
    + tnln=0.06811233782202991u tnwn=112.0090347746391n tnotv=1.6768540479291394n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.07246753667703952u tpotv=1.7845041168722293n tpwv=226.76492451036412n 
    + tnln=0.06523301181742534u tnwn=130.41129396195603n tnotv=1.9793945985792736n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.07389910284973608u tpotv=1.8834224689870749n tpwv=200.4725084365421n 
    + tnln=0.05563790034761337u tnwn=122.06325122519394n tnotv=2.0203730008200877n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06317983543191742u tpotv=2.011916708122805n tpwv=236.40717387261847n 
    + tnln=0.05915969422410062u tnwn=128.29436794432777n tnotv=1.850908380715777n 

.ENDS ring_osc.end
