* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_0 in0 out12 vdd 0

    x0 in0 out12 out0 vdd 0 nand params:
    + tplv=0.06716981076063507u tpotv=2.1359217630130294n tpwv=119.76360958021269n 
    + tnln=0.06913924322856611u tnwn=123.44118827616566n tnotv=1.9370273403402898n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.07132370359557018u tpotv=2.0649526300647816n tpwv=243.10821640449643n 
    + tnln=0.07331727464256388u tnwn=136.15558883167193n tnotv=1.8408663108688743n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.055882264060639335u tpotv=1.8673884657752882n tpwv=248.10014142775995n 
    + tnln=0.0612270663088998u tnwn=141.40104575975235n tnotv=1.841415275228472n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06111244788915603u tpotv=2.0264757055189553n tpwv=186.13262302341593n 
    + tnln=0.06525650413595463u tnwn=142.9705636533821n tnotv=1.946333197418418n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.06800359808431763u tpotv=1.8422740836365428n tpwv=206.99062393715474n 
    + tnln=0.06604057260806286u tnwn=117.94431913153765n tnotv=1.9447755643302231n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.07374839555060672u tpotv=1.8111185593704209n tpwv=205.35928544286676n 
    + tnln=0.0728127023566856u tnwn=129.41862977928184n tnotv=1.6684214369450838n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.05860597651325626u tpotv=1.8726136995609195n tpwv=248.90855337236786n 
    + tnln=0.060712252979839024u tnwn=121.44334413738534n tnotv=2.021738423177273n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.07116305078202813u tpotv=2.138345629994694n tpwv=205.35794117948114n 
    + tnln=0.0740538912159624u tnwn=139.34085266297248n tnotv=2.018914011408474n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.0684449302946091u tpotv=2.021682562582617n tpwv=190.8174566743511n 
    + tnln=0.056825614538021485u tnwn=127.99451683101631n tnotv=1.7554587077790909n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0665482941725159u tpotv=1.9269915183827864n tpwv=207.8581062732135n 
    + tnln=0.05689187546830611u tnwn=115.8673254150179n tnotv=1.9702843711186868n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06735634268634007u tpotv=1.9564132385001536n tpwv=208.98673670936176n 
    + tnln=0.07471361193658778u tnwn=121.69876855775772n tnotv=1.7784741398069972n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.06733617134181187u tpotv=1.9402441779987503n tpwv=241.34449768025829n 
    + tnln=0.05587662495988516u tnwn=130.37391695363397n tnotv=1.9592275834419177n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.05633887325674055u tpotv=1.8650690244300312n tpwv=186.96378200862398n 
    + tnln=0.05570275211041394u tnwn=131.36180492259925n tnotv=1.7309921327209814n 

.ENDS ring_osc.end
