* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_0 in0 out12 vdd 0

    x0 in0 out12 out0 vdd 0 nand params:
    + tplv=0.06767110151070026u tpotv=1.8005034378768916n tpwv=114.38439228295617n 
    + tnln=0.0686369587980066u tnwn=116.65287488874537n tnotv=1.8354339464191851n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.0557934964539917u tpotv=1.8433717610980214n tpwv=187.65866748605657n 
    + tnln=0.06979895696959312u tnwn=147.70500295423142n tnotv=1.9612456836015342n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06738434262077352u tpotv=2.0086975785552466n tpwv=211.47237767101782n 
    + tnln=0.0676658227519368u tnwn=142.2660332722838n tnotv=1.6958194380691447n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.05922518763974732u tpotv=1.9840064289716555n tpwv=244.6056493308454n 
    + tnln=0.05950229790993298u tnwn=133.06705663634068n tnotv=1.9390360641085407n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.05921108879605054u tpotv=1.9741544819859624n tpwv=188.95987679738187n 
    + tnln=0.05722929154681344u tnwn=131.48482006702355n tnotv=1.678683253759526n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.072105084157307u tpotv=1.9225785007772065n tpwv=191.16238805076222n 
    + tnln=0.06018602298251727u tnwn=133.88255146700672n tnotv=1.7799682228497336n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.0674145290723994u tpotv=2.082330053075003n tpwv=194.38714396129967n 
    + tnln=0.05801103520286188u tnwn=133.76779397633396n tnotv=1.713003681762203n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.07261179703521706u tpotv=2.070087806287021n tpwv=228.45058152802238n 
    + tnln=0.07293561505480368u tnwn=127.58000184902205n tnotv=1.962892806143291n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.062465090853928554u tpotv=1.8375485372433134n tpwv=195.76392598547685n 
    + tnln=0.06245961165697925u tnwn=123.62811074459219n tnotv=1.7480286698282734n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06067305596429101u tpotv=1.9171662931534275n tpwv=229.22102147062913n 
    + tnln=0.0649689960806831u tnwn=143.05713309128996n tnotv=1.7721525088204468n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06805782749213048u tpotv=1.8418850355550307n tpwv=232.7672774841221n 
    + tnln=0.06933469193131843u tnwn=124.58631745749992n tnotv=1.945665504550762n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.06443315154833273u tpotv=1.9768052713286917n tpwv=188.9028517558985n 
    + tnln=0.058994254151581646u tnwn=115.77386180777845n tnotv=1.7335948756073258n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.05740926491227126u tpotv=1.9539481588690284n tpwv=205.21493364376676n 
    + tnln=0.06300741039986782u tnwn=148.13666346235146n tnotv=1.9949886230867597n 

.ENDS ring_osc.end
