* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_1 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.07173908243594779u tpotv=1.826112067640427n tpwv=250.08595093623066n 
    + tnln=0.06502695278571594u tnwn=123.17321542814992n tnotv=1.9112180092546145n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.07323722561860838u tpotv=2.1020060351065823n tpwv=217.77305892884684n 
    + tnln=0.06562323440231627u tnwn=121.75745280130232n tnotv=1.776906323850783n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.07416286451579286u tpotv=1.853315155558239n tpwv=248.2000905375031n 
    + tnln=0.06727624266412616u tnwn=119.8191431229367n tnotv=1.8387866220792812n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.061847191327190694u tpotv=2.057384992488828n tpwv=198.5630013210978n 
    + tnln=0.05562593579483684u tnwn=134.96611155760615n tnotv=2.0198906521314774n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.057460663821183415u tpotv=2.034257216226606n tpwv=230.2445115979319n 
    + tnln=0.05842180608030528u tnwn=111.71317462618987n tnotv=1.8168021001485386n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06193049064177827u tpotv=1.800519849454819n tpwv=241.82147844271708n 
    + tnln=0.06834121982431057u tnwn=121.74336974673372n tnotv=1.9034380718524586n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06059141289094276u tpotv=1.9630388985128167n tpwv=211.50426612412713n 
    + tnln=0.06730879535504926u tnwn=135.5926823864637n tnotv=1.7311725624150083n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06778214439881233u tpotv=1.9296319209140536n tpwv=220.41404538609066n 
    + tnln=0.06829931963446968u tnwn=110.6228579782591n tnotv=1.7727068744874364n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.07347015360526332u tpotv=2.0368975711786974n tpwv=193.61130859333747n 
    + tnln=0.06018218737854575u tnwn=116.35382611668652n tnotv=2.024878672872333n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0700824231708684u tpotv=2.0806886887930065n tpwv=246.79891552884888n 
    + tnln=0.055591657615030404u tnwn=130.12018615940516n tnotv=1.9611037464347296n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.07413476475346541u tpotv=2.0097805393373047n tpwv=248.91521820293855n 
    + tnln=0.06344799124805978u tnwn=132.96265483757745n tnotv=2.0115673702910093n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.05900331267453124u tpotv=1.948406424285706n tpwv=221.9182916706103n 
    + tnln=0.07413997546696553u tnwn=133.67579016174506n tnotv=1.9995276303925746n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.07355806727229493u tpotv=1.8330842661167788n tpwv=237.52962552981174n 
    + tnln=0.0708289854195348u tnwn=125.56456076673217n tnotv=1.974482234687937n 

.ENDS ring_osc.end
