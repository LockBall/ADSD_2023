
module TSD_ADC (
	clk_clk,
	reset_reset_n,
	altpll_0_inclk_interface_clk,
	altpll_0_inclk_interface_reset_reset);	

	input		clk_clk;
	input		reset_reset_n;
	input		altpll_0_inclk_interface_clk;
	input		altpll_0_inclk_interface_reset_reset;
endmodule
