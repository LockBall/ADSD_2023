* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_7 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.06818285569813819u tpotv=2.0306291589512573n tpwv=226.7654419310441n 
    + tnln=0.06167128041016384u tnwn=115.48821103929568n tnotv=2.0110913294960646n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06885145926821681u tpotv=2.0023431027283998n tpwv=225.52305692284733n 
    + tnln=0.07410362093657007u tnwn=134.76401537116857n tnotv=1.684549259767173n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.05588585785299745u tpotv=1.828497006833752n tpwv=232.85682394092984n 
    + tnln=0.06505548643279792u tnwn=137.7064091504812n tnotv=1.9631686782603053n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.07377081822758257u tpotv=1.8647612216993865n tpwv=219.4175814366965n 
    + tnln=0.07213325698886691u tnwn=138.04609723371252n tnotv=1.900170709258808n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.07280519508842703u tpotv=1.8715731604388848n tpwv=231.48633750694893n 
    + tnln=0.06720465869431323u tnwn=141.5406726789519n tnotv=2.0317139723048525n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.07235191520620331u tpotv=1.8493882715749954n tpwv=227.95865132389733n 
    + tnln=0.05892144472121927u tnwn=118.80010155088013n tnotv=1.6982315373109373n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.057442548667872184u tpotv=1.9172875137703966n tpwv=246.92308607918426n 
    + tnln=0.0739267639752957u tnwn=123.9670073537245n tnotv=1.7246396930746026n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06032556019813017u tpotv=1.8720781797549417n tpwv=249.65304470583166n 
    + tnln=0.0581319563585124u tnwn=145.0027654884356n tnotv=1.6842661137060815n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06781049571888882u tpotv=2.122406249212498n tpwv=230.64501894846154n 
    + tnln=0.06477006489034617u tnwn=113.83899715621915n tnotv=1.755342607887445n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.0736640734186954u tpotv=2.0135596359773253n tpwv=211.5333412240551n 
    + tnln=0.06687150685196826u tnwn=136.9228215698996n tnotv=1.9007431012086198n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.05847411329114257u tpotv=2.1374766323091876n tpwv=185.87027197913514n 
    + tnln=0.05698797203000845u tnwn=111.36927784057158n tnotv=1.7068647179249146n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.07279759123038722u tpotv=1.934104125527805n tpwv=203.85767193761336n 
    + tnln=0.061692473387221114u tnwn=118.41678326698215n tnotv=1.846755676538621n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06834236325901848u tpotv=1.8937163909002512n tpwv=210.2607671886929n 
    + tnln=0.06683001005902847u tnwn=136.88758275553914n tnotv=1.7539554486755062n 

.ENDS ring_osc.end
