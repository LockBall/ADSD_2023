* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_6 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.06716308410975741u tpotv=2.0969308930963737n tpwv=230.76030546706684n 
    + tnln=0.06432662891994528u tnwn=131.4346527142232n tnotv=1.852971324887075n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06820273592280596u tpotv=1.9365524904016858n tpwv=200.52418011134822n 
    + tnln=0.07128322450032212u tnwn=126.27362162427323n tnotv=1.82217636562644n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.05638073171273501u tpotv=1.7632119442276215n tpwv=196.6138655227916n 
    + tnln=0.062005198453554185u tnwn=129.54831406051883n tnotv=1.6902084311403487n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.07276956031000935u tpotv=1.8808430376529437n tpwv=198.08976265023767n 
    + tnln=0.07178958266121821u tnwn=135.11097967637323n tnotv=1.697073376770256n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.06591005964068887u tpotv=1.895085813967908n tpwv=226.0263525212434n 
    + tnln=0.05699610584533321u tnwn=123.59712130193584n tnotv=1.9340029852594913n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.0729069091912048u tpotv=1.8991409574233846n tpwv=234.10851397766038n 
    + tnln=0.05719538575319327u tnwn=125.51308276474577n tnotv=1.8084853538335672n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06841602896157072u tpotv=2.0877472984602643n tpwv=228.8295818431313n 
    + tnln=0.06355110559850623u tnwn=140.17808931310512n tnotv=2.0174648374976614n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.059177533847321225u tpotv=1.8131433980614666n tpwv=234.5263753292722n 
    + tnln=0.06006625103941472u tnwn=141.71862203843654n tnotv=2.0248371898985575n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06528134528174166u tpotv=2.0929155057694775n tpwv=239.23790354722505n 
    + tnln=0.06704161961557949u tnwn=134.2311020543975n tnotv=1.891395458875285n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.07188681615082032u tpotv=1.9316257009467541n tpwv=229.11826254119225n 
    + tnln=0.0580980130919385u tnwn=130.22987464926837n tnotv=2.009589378642827n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.05994538478188228u tpotv=1.9436770314636869n tpwv=194.9652774642497n 
    + tnln=0.06374622987272736u tnwn=130.42447294137n tnotv=1.6750439594645479n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.0641084275147595u tpotv=2.0385774595698836n tpwv=214.40495818341574n 
    + tnln=0.058018752185897485u tnwn=142.6823388454602n tnotv=1.8659385759120426n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.07417304483924995u tpotv=1.8356239679175848n tpwv=243.77970231792688n 
    + tnln=0.06394988293042854u tnwn=129.57675204211594n tnotv=1.8165753636670021n 

.ENDS ring_osc.end
