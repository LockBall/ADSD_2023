clock_10_inst : clock_10 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
