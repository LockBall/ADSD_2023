* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_5 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.061028903045290836u tpotv=1.7687484962870788n tpwv=246.7244837439096n 
    + tnln=0.05722267534996413u tnwn=111.82621578539272n tnotv=1.6800147825172038n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.0681904332112005u tpotv=1.8670879836695826n tpwv=237.08816650310817n 
    + tnln=0.07156619403404119u tnwn=147.31733407767865n tnotv=1.9279240680315222n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06405739633930785u tpotv=1.9476143529477332n tpwv=216.28191804760866n 
    + tnln=0.06016033232677136u tnwn=112.8831317722769n tnotv=1.7487237319437348n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.056538078493041245u tpotv=1.8619355722524695n tpwv=232.459660224476n 
    + tnln=0.07086400171179845u tnwn=110.64278389361735n tnotv=1.842722791361014n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.058199738453835026u tpotv=2.082786798184286n tpwv=211.908524879358n 
    + tnln=0.06681622874757592u tnwn=134.77742051192257n tnotv=1.793993126530648n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.07058615173927679u tpotv=1.9603286514673721n tpwv=235.38616294659224n 
    + tnln=0.05984694462330095u tnwn=138.80597083675033n tnotv=1.696561828028943n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.05615282495384917u tpotv=1.898248019947467n tpwv=220.2742123120993n 
    + tnln=0.058744076647988405u tnwn=117.97631954647528n tnotv=1.896885859335895n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.05918152605466198u tpotv=1.7717764265018947n tpwv=207.87047374410338n 
    + tnln=0.07025937941389047u tnwn=130.28192957706233n tnotv=1.9627129568919628n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06751053808942664u tpotv=1.9363047387050665n tpwv=215.20571601819577n 
    + tnln=0.06051665285772313u tnwn=139.765814601803n tnotv=1.9635642301098921n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06417398358483245u tpotv=2.0520941645120727n tpwv=189.37468081969342n 
    + tnln=0.06076278319944603u tnwn=139.09575910538265n tnotv=1.8256386720942919n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06531112552239034u tpotv=2.0668624303326877n tpwv=207.39836809309043n 
    + tnln=0.055352100367245236u tnwn=121.40379432769069n tnotv=1.8870781675597408n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.061887584626078504u tpotv=1.7805329203563476n tpwv=190.47107784570198n 
    + tnln=0.056742817774847104u tnwn=141.70965597372881n tnotv=1.9207889390423885n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06168758639955574u tpotv=1.7644845269533875n tpwv=237.31463056263763n 
    + tnln=0.06259932845615562u tnwn=111.66048308978463n tnotv=1.7128412304881657n 

.ENDS ring_osc.end
