* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_4 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.07429581688222128u tpotv=1.8375229060243856n tpwv=225.4003550938359n 
    + tnln=0.056911110290462745u tnwn=145.86217819698587n tnotv=1.964040751579441n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06278979077279362u tpotv=2.090399354802407n tpwv=225.56322643047872n 
    + tnln=0.05908228975301237u tnwn=127.87583621748976n tnotv=2.0267487166001046n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.05659842725345712u tpotv=2.021300430482991n tpwv=218.96128666496716n 
    + tnln=0.05558840586137055u tnwn=133.75633733905076n tnotv=2.0174474772796267n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06434676081185839u tpotv=2.0011066673266584n tpwv=209.76619981247734n 
    + tnln=0.05932657852637298u tnwn=131.85952162171523n tnotv=1.7299829160779885n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.05572822823960372u tpotv=1.7659402095292478n tpwv=243.72324370042924n 
    + tnln=0.06838457093853824u tnwn=122.43661804948576n tnotv=2.0061342106259237n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.05746907247468411u tpotv=1.8661289358757511n tpwv=248.8775374123732n 
    + tnln=0.06514050820283154u tnwn=147.90716048240634n tnotv=1.9665236478653072n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.05642408678419811u tpotv=1.8473637915006536n tpwv=223.11399565106615n 
    + tnln=0.06404819570614466u tnwn=143.04464193040394n tnotv=1.9957937406857942n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.055603432826809546u tpotv=2.130443461744703n tpwv=198.54445658481052n 
    + tnln=0.06190246293618148u tnwn=118.69707271716092n tnotv=2.0044423261163695n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.057382524718292194u tpotv=1.908118989170658n tpwv=226.35570142425752n 
    + tnln=0.07025371031390461u tnwn=148.19776328107898n tnotv=1.8427089002206385n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.07209162625969061u tpotv=1.931008064883416n tpwv=196.2992329453762n 
    + tnln=0.07401875711418648u tnwn=117.65594588954113n tnotv=1.775314384104593n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.07207945200076263u tpotv=2.1389392776366822n tpwv=207.7484015197011n 
    + tnln=0.06881958033818822u tnwn=111.83724030288724n tnotv=1.8242205231557975n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.057790044615729994u tpotv=1.8486270083084477n tpwv=218.34802810277205n 
    + tnln=0.056201017082906944u tnwn=137.51010012881378n tnotv=1.9381314902520361n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.07127056982199241u tpotv=2.1115213083427n tpwv=203.73815411480723n 
    + tnln=0.07138699836416736u tnwn=148.0034089195401n tnotv=1.984687346596934n 

.ENDS ring_osc.end
