* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_7 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.0698056323007993u tpotv=2.0023256791657085n tpwv=217.39503277489n 
    + tnln=0.06504316354215435u tnwn=144.5075341795125n tnotv=1.8915947412628245n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06013955882266403u tpotv=1.8254945986465092n tpwv=217.13758446336178n 
    + tnln=0.06546717676835798u tnwn=147.27234545674312n tnotv=1.8642636864549986n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.0743122989401612u tpotv=1.9345368238548777n tpwv=186.62212145313313n 
    + tnln=0.056133743109334146u tnwn=115.90851010873038n tnotv=1.8182125373320106n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.05556033515542593u tpotv=2.022072293192794n tpwv=202.15384183544398n 
    + tnln=0.06703816526449148u tnwn=116.72060734238329n tnotv=1.963964659168931n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.07200140017074069u tpotv=1.8843839547323606n tpwv=215.09272977455817n 
    + tnln=0.07368482286612406u tnwn=112.8253861241274n tnotv=1.9735499556874507n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06338400984096446u tpotv=1.9246178499932611n tpwv=219.58477392636416n 
    + tnln=0.07386113105289803u tnwn=112.3363984757699n tnotv=1.7381639912134954n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06258794215575489u tpotv=2.085573615943717n tpwv=230.06130661589756n 
    + tnln=0.06323099330864042u tnwn=131.49646783805636n tnotv=1.6809837551316167n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06074030929960203u tpotv=1.8073711741159588n tpwv=242.6882255181878n 
    + tnln=0.06976152817480397u tnwn=148.63382570067887n tnotv=1.6662989546850873n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.06930150457985557u tpotv=1.7558706783854348n tpwv=237.328144079948n 
    + tnln=0.06443674847101763u tnwn=111.43719186192133n tnotv=1.8582898087121502n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06752238065087457u tpotv=1.9260723359562224n tpwv=247.188543461628n 
    + tnln=0.06531591650385435u tnwn=111.11824205548965n tnotv=1.9962080321631241n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.07047972756928868u tpotv=1.944169976003038n tpwv=227.8038186372296n 
    + tnln=0.06158914153322209u tnwn=128.7069912394884n tnotv=1.7386916260977796n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.06630111252498404u tpotv=1.8463101971673206n tpwv=241.74410085381726n 
    + tnln=0.07200697612574669u tnwn=141.89539800065847n tnotv=1.9545760213046837n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.061282713228595895u tpotv=1.9955975464866258n tpwv=241.62239181706553n 
    + tnln=0.07329272459428235u tnwn=125.20190056705536n tnotv=1.9291055739239051n 

.ENDS ring_osc.end
