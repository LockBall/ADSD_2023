* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_2 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.06287967379300159u tpotv=2.016640610822183n tpwv=232.7666924825977n 
    + tnln=0.06124716321447141u tnwn=126.34394437937591n tnotv=1.6794379795885268n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06696141905984387u tpotv=2.047684904247913n tpwv=237.37500970468366n 
    + tnln=0.07403283507004821u tnwn=115.4515690783604n tnotv=1.8734481997415082n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.05857571165943133u tpotv=2.0038126076970912n tpwv=202.59484936107464n 
    + tnln=0.0676001550378642u tnwn=144.46354037921571n tnotv=1.9947551366089828n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.05997073430801833u tpotv=1.9507437522827122n tpwv=217.47754211342547n 
    + tnln=0.06657767184369552u tnwn=119.56823288139269n tnotv=1.735068766564619n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.0662222723259539u tpotv=1.9006409292455144n tpwv=214.57619260434885n 
    + tnln=0.06798538818634486u tnwn=116.32914076213402n tnotv=1.964898649221185n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.07048898690617679u tpotv=2.1194395982940293n tpwv=187.45545127417876n 
    + tnln=0.05607920629244155u tnwn=141.5061912160062n tnotv=1.6697797668214953n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.06792177584163092u tpotv=2.066326187299364n tpwv=226.27821569400822n 
    + tnln=0.061182599009036984u tnwn=135.98310073052855n tnotv=1.806185926961179n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.06716057451477325u tpotv=2.1042153114534785n tpwv=225.57203263164604n 
    + tnln=0.061064600243168565u tnwn=147.18162780955407n tnotv=1.898421388656729n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.062184885474295216u tpotv=1.8428416896348938n tpwv=219.6735689222596n 
    + tnln=0.0573977945528069u tnwn=122.87010972261339n tnotv=1.7460207543789248n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.06551441447561789u tpotv=2.0746184846452254n tpwv=232.55486295784866n 
    + tnln=0.07075834687277145u tnwn=120.93037044688649n tnotv=1.9352318729608848n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06862703129267757u tpotv=1.9601114707150766n tpwv=193.03679373085805n 
    + tnln=0.06342191279570118u tnwn=131.7082055936922n tnotv=1.9007567582748057n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.0674897165534249u tpotv=1.8939336929222939n tpwv=189.65344692604688n 
    + tnln=0.06523359691478409u tnwn=137.69526339238467n tnotv=1.6690288174277006n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06324859890200646u tpotv=1.8426553049679364n tpwv=235.18551375254373n 
    + tnln=0.06564834975712898u tnwn=139.7120201086035n tnotv=1.7405132426033214n 

.ENDS ring_osc.end
