library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;


library floatfixlib;
use floatfixlib.fixed_pkg.all;

entity mando_ppm is



architecture arch of mando_ppm is

-- signals

  begin
  
  

end arch ;