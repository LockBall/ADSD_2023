* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_3 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.060314261989083615u tpotv=1.9213556872399173n tpwv=236.61942701973086n 
    + tnln=0.06597573096865614u tnwn=119.98516244755274n tnotv=1.748907258051696n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.06205911572686342u tpotv=1.7670750909749589n tpwv=190.02346765866582n 
    + tnln=0.06743472635549744u tnwn=127.29378074242386n tnotv=1.7122175783962157n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.06565975570956323u tpotv=2.0532687479510225n tpwv=233.98506680103634n 
    + tnln=0.056653133701339634u tnwn=144.48721055253478n tnotv=1.9117965405261916n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06492993517795874u tpotv=1.891769294536238n tpwv=194.0684132224231n 
    + tnln=0.06191668412140523u tnwn=142.99831673569562n tnotv=1.6743498855858248n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.06887273014146844u tpotv=2.0424032869513216n tpwv=219.4571790056383n 
    + tnln=0.05637857399160777u tnwn=111.1829447215849n tnotv=1.978609122743964n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06073493942918723u tpotv=1.7899992370404303n tpwv=193.74549197066085n 
    + tnln=0.060913701335227784u tnwn=116.45269289768227n tnotv=1.7003595199992885n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.0601180597451336u tpotv=1.7697981652936257n tpwv=214.58526305331048n 
    + tnln=0.06573709242819534u tnwn=134.10130346076662n tnotv=1.9518778268220773n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.05943963516465574u tpotv=2.072148236280387n tpwv=221.8035510565771n 
    + tnln=0.06750934890741332u tnwn=130.37309350947157n tnotv=1.862014225771381n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.060988840493991024u tpotv=2.0833047705681658n tpwv=200.39037973361863n 
    + tnln=0.07196777439990454u tnwn=140.83385185501507n tnotv=1.6783895838295426n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.05560511898756523u tpotv=1.950855652673411n tpwv=218.06370939071226n 
    + tnln=0.07451142053485216u tnwn=125.64696757917241n tnotv=1.924761369946779n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.06398659384178283u tpotv=2.0946291371627597n tpwv=188.87240769865858n 
    + tnln=0.07116096974873705u tnwn=127.54924200183345n tnotv=1.8035460063723183n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.06904802182606917u tpotv=2.1185464775873544n tpwv=249.69557443006417n 
    + tnln=0.06589398912654522u tnwn=135.39962649905937n tnotv=1.6770037656327965n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.07470225721906963u tpotv=1.8770501452078074n tpwv=244.5175575719923n 
    + tnln=0.0562923589406351u tnwn=144.6250159299005n tnotv=1.7817733858881315n 

.ENDS ring_osc.end
