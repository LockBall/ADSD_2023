* Generator created 01 Oct 2022 by John Lutz. Editeded 02 Oct 2022
* This file generated on: 13 Sep 2023

.SUBCKT ring_osc_5 in0 out12 vdd 0

    x0 in0 out0 vdd 0 inverter params:
    + tplv=0.07443550772050495u tpotv=1.806151139931906n tpwv=241.2635436559237n 
    + tnln=0.05842430377447576u tnwn=118.08390814749997n tnotv=1.9606529746893282n 

    x1 out0 out1 vdd 0 inverter params:
    + tplv=0.0650970572479821u tpotv=1.8168741116643652n tpwv=216.47178211355563n 
    + tnln=0.059984416667260176u tnwn=142.26875119150557n tnotv=2.012069560159998n 

    x2 out1 out2 vdd 0 inverter params:
    + tplv=0.0632944521462687u tpotv=2.1107045995494955n tpwv=216.61792646536944n 
    + tnln=0.056717938845173684u tnwn=122.41658961914027n tnotv=1.731287776964738n 

    x3 out2 out3 vdd 0 inverter params:
    + tplv=0.06433111145549178u tpotv=2.1224299413339462n tpwv=231.48783118816417n 
    + tnln=0.07259299292180865u tnwn=117.89733643303475n tnotv=1.914245094177832n 

    x4 out3 out4 vdd 0 inverter params:
    + tplv=0.05532945973470789u tpotv=2.032480680011984n tpwv=224.694256532145n 
    + tnln=0.0743255800520983u tnwn=119.29467468772863n tnotv=1.7698331973773944n 

    x5 out4 out5 vdd 0 inverter params:
    + tplv=0.06517202802281132u tpotv=1.9799296270638334n tpwv=242.0468792648131n 
    + tnln=0.06435385403788119u tnwn=139.87877783601186n tnotv=2.016621143265951n 

    x6 out5 out6 vdd 0 inverter params:
    + tplv=0.07324018865161326u tpotv=1.9807626389587862n tpwv=217.51837403451054n 
    + tnln=0.07242367023642315u tnwn=146.8573112785588n tnotv=1.9401056897457882n 

    x7 out6 out7 vdd 0 inverter params:
    + tplv=0.0593357306669291u tpotv=1.7823340055239714n tpwv=247.71440134574092n 
    + tnln=0.07078564448538271u tnwn=147.24031075774306n tnotv=1.9480372343554617n 

    x8 out7 out8 vdd 0 inverter params:
    + tplv=0.05739908580993883u tpotv=2.112246729681981n tpwv=216.8956902425743n 
    + tnln=0.07442820606034356u tnwn=127.9133992871943n tnotv=1.756973632586606n 

    x9 out8 out9 vdd 0 inverter params:
    + tplv=0.05831766515343761u tpotv=2.06190263680212n tpwv=211.27266085514952n 
    + tnln=0.05852478638295927u tnwn=137.76845312451584n tnotv=1.9868968693558269n 

    x10 out9 out10 vdd 0 inverter params:
    + tplv=0.057177155757345284u tpotv=2.0314432315405755n tpwv=193.51892908219202n 
    + tnln=0.07204992859699337u tnwn=123.82371490711489n tnotv=1.9991205615148155n 

    x11 out10 out11 vdd 0 inverter params:
    + tplv=0.07246934471660336u tpotv=1.9064406105112135n tpwv=236.55594437590707n 
    + tnln=0.05842760263653772u tnwn=116.41339665354721n tnotv=1.9239937888778103n 

    x12 out11 out12 vdd 0 inverter params:
    + tplv=0.06457465922291951u tpotv=1.782366260559548n tpwv=187.5736303731487n 
    + tnln=0.055772997180055406u tnwn=124.54459560317198n tnotv=1.998260556944491n 

.ENDS ring_osc.end
